module alu_simple_tb;

    // ====================================================================
    // ส่วนที่ 1: ประกาศสัญญาณ
    // ====================================================================
    // ✅ ถูกต้องแล้ว!
    reg  [31:0] A;
    reg  [31:0] B;
    reg  [1:0]  ALUControl;
    wire [31:0] Result;
    wire        Zero;

    // ====================================================================
    // ส่วนที่ 2: Instance ของ ALU
    // ====================================================================
    // ✅ ดีมาก! ชื่อ dut (Design Under Test) เป็นมาตรฐาน
    alu_simple dut (
        .A(A),
        .B(B),
        .ALUControl(ALUControl),
        .Result(Result),
        .Zero(Zero)
    );

    // ====================================================================
    // ส่วนที่ 3: Monitor
    // ====================================================================
    // ✅ ดี! แต่ปรับปรุงให้อ่านง่ายขึ้น
    initial begin
        $display("=================================================================");
        $display("🧪 เริ่มทดสอบ ALU");
        $display("=================================================================");
        $display("Time | Control | Operation |    A    |    B    |  Result | Zero");
        $display("-----------------------------------------------------------------");
    end
    
    // Monitor แสดงผลทุกครั้งที่มีการเปลี่ยนแปลง
    always @(A, B, ALUControl, Result, Zero) begin
        // หน่วงเวลาเล็กน้อยเพื่อให้ผลลัพธ์เสถียร
        #1;
        
        // แสดงชื่อ operation ให้เข้าใจง่าย
        case(ALUControl)
            2'b00: $display("%4t |   %b    |    AND    | %7d | %7d | %7d |  %b",
                           $time, ALUControl, A, B, Result, Zero);
            2'b01: $display("%4t |   %b    |    OR     | %7d | %7d | %7d |  %b",
                           $time, ALUControl, A, B, Result, Zero);
            2'b10: $display("%4t |   %b    |    ADD    | %7d | %7d | %7d |  %b",
                           $time, ALUControl, A, B, Result, Zero);
            2'b11: $display("%4t |   %b    |    SUB    | %7d | %7d | %7d |  %b",
                           $time, ALUControl, A, B, Result, Zero);
        endcase
    end

    // ====================================================================
    // ส่วนที่ 4: Test Vectors
    // ====================================================================
    initial begin
        // เริ่มต้นค่า
        A = 32'd0;
        B = 32'd0;
        ALUControl = 2'b00;
        
        // --------------------------------------------------------
        // Test 1: AND
        // --------------------------------------------------------
        #10;
        $display("\n--- Test 1: AND ---");
        A = 32'd10;         // 0000...1010
        B = 32'd5;          // 0000...0101
        ALUControl = 2'b00; // AND
        #10;
        $display("คำอธิบาย: 1010 & 0101 = 0000 (ทศนิยม = 0)");
        
        // --------------------------------------------------------
        // Test 2: OR
        // --------------------------------------------------------
        $display("\n--- Test 2: OR ---");
        A = 32'd10;         // 0000...1010
        B = 32'd5;          // 0000...0101
        ALUControl = 2'b01; // OR
        #10;
        $display("คำอธิบาย: 1010 | 0101 = 1111 (ทศนิยม = 15)");
        
        // --------------------------------------------------------
        // Test 3: ADD
        // --------------------------------------------------------
        $display("\n--- Test 3: ADD ---");
        A = 32'd10;
        B = 32'd5;
        ALUControl = 2'b10; // ADD
        #10;
        $display("คำอธิบาย: 10 + 5 = 15 ✅");
        
        // --------------------------------------------------------
        // Test 4: SUB
        // --------------------------------------------------------
        $display("\n--- Test 4: SUB ---");
        A = 32'd10;
        B = 32'd5;
        ALUControl = 2'b11; // SUB
        #10;
        $display("คำอธิบาย: 10 - 5 = 5 ✅");
        
        // --------------------------------------------------------
        // Test 5: Zero Flag (ผลลัพธ์เป็นศูนย์)
        // --------------------------------------------------------
        $display("\n--- Test 5: SUB → Zero Flag ---");
        A = 32'd8;
        B = 32'd8;
        ALUControl = 2'b11; // SUB
        #10;
        $display("คำอธิบาย: 8 - 8 = 0 → Zero = 1 ✅");
        
        // --------------------------------------------------------
        // Test 6: ผลลัพธ์ติดลบ
        // --------------------------------------------------------
        $display("\n--- Test 6: SUB → Negative Result ---");
        A = 32'd5;
        B = 32'd10;
        ALUControl = 2'b11; // SUB
        #10;
        $display("คำอธิบาย: 5 - 10 = -5");
        $display("ในระบบ 2's complement: Result = %d", $signed(Result));
        
        // --------------------------------------------------------
        // Test 7: เลขใหญ่
        // --------------------------------------------------------
        $display("\n--- Test 7: ADD → Large Numbers ---");
        A = 32'd1000000;
        B = 32'd2000000;
        ALUControl = 2'b10; // ADD
        #10;
        $display("คำอธิบาย: 1,000,000 + 2,000,000 = 3,000,000 ✅");
        
        // --------------------------------------------------------
        // จบการทดสอบ
        // --------------------------------------------------------
        #10;
        $display("\n=================================================================");
        $display("🎉 ทดสอบเสร็จสมบูรณ์!");
        $display("=================================================================");
        $display("\n📊 สรุป:");
        $display("   ✅ AND  - ทดสอบแล้ว");
        $display("   ✅ OR   - ทดสอบแล้ว");
        $display("   ✅ ADD  - ทดสอบแล้ว");
        $display("   ✅ SUB  - ทดสอบแล้ว");
        $display("   ✅ Zero Flag - ทดสอบแล้ว");
        $display("   ✅ Negative - ทดสอบแล้ว");
        $display("\n");
        
        $finish;
    end

endmodule